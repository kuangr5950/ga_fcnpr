module c432 ( 
    \1 , 4, 8, 11, 14, 17, 21, 24, 27, 30, 34, 37, 40, 43, 47, 50, 53, 56,
    60, 63, 66, 69, 73, 76, 79, 82, 86, 89, 92, 95, 99, 102, 105, 108, 112,
    115,
    223, 329, 370, 421, 430, 431, 432  );
  input  \1 , 4, 8, 11, 14, 17, 21, 24, 27, 30, 34, 37, 40, 43, 47, 50,
    53, 56, 60, 63, 66, 69, 73, 76, 79, 82, 86, 89, 92, 95, 99, 102, 105,
    108, 112, 115;
  output 223, 329, 370, 421, 430, 431, 432;
  wire n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
    n58, n59, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n238, n239, n241, n242, n243, n244, n245, n246, n248, n249,
    n250, n251;
  assign n44 = ~\1  & 4;
  assign n45 = ~11 & 17;
  assign n46 = ~24 & 30;
  assign n47 = ~37 & 43;
  assign n48 = ~50 & 56;
  assign n49 = ~63 & 69;
  assign n50 = ~76 & 82;
  assign n51 = ~89 & 95;
  assign n52 = ~102 & 108;
  assign n53 = ~n44 & ~n45;
  assign n54 = ~n46 & n53;
  assign n55 = ~n47 & n54;
  assign n56 = ~n48 & n55;
  assign n57 = ~n49 & n56;
  assign n58 = ~n50 & n57;
  assign n59 = ~n51 & n58;
  assign 223 = n52 | ~n59;
  assign n61 = ~n44 & ~223;
  assign n62 = n44 & 223;
  assign n63 = ~n61 & ~n62;
  assign n64 = 4 & ~8;
  assign n65 = ~n63 & n64;
  assign n66 = ~n45 & ~223;
  assign n67 = n45 & 223;
  assign n68 = ~n66 & ~n67;
  assign n69 = 17 & ~21;
  assign n70 = ~n68 & n69;
  assign n71 = ~n46 & ~223;
  assign n72 = n46 & 223;
  assign n73 = ~n71 & ~n72;
  assign n74 = 30 & ~34;
  assign n75 = ~n73 & n74;
  assign n76 = ~n47 & ~223;
  assign n77 = n47 & 223;
  assign n78 = ~n76 & ~n77;
  assign n79 = 43 & ~47;
  assign n80 = ~n78 & n79;
  assign n81 = ~n48 & ~223;
  assign n82 = n48 & 223;
  assign n83 = ~n81 & ~n82;
  assign n84 = 56 & ~60;
  assign n85 = ~n83 & n84;
  assign n86 = ~n49 & ~223;
  assign n87 = n49 & 223;
  assign n88 = ~n86 & ~n87;
  assign n89 = 69 & ~73;
  assign n90 = ~n88 & n89;
  assign n91 = ~n50 & ~223;
  assign n92 = n50 & 223;
  assign n93 = ~n91 & ~n92;
  assign n94 = 82 & ~86;
  assign n95 = ~n93 & n94;
  assign n96 = ~n51 & ~223;
  assign n97 = n51 & 223;
  assign n98 = ~n96 & ~n97;
  assign n99 = 95 & ~99;
  assign n100 = ~n98 & n99;
  assign n101 = ~n52 & ~223;
  assign n102 = n52 & 223;
  assign n103 = ~n101 & ~n102;
  assign n104 = 108 & ~112;
  assign n105 = ~n103 & n104;
  assign n106 = ~n65 & ~n70;
  assign n107 = ~n75 & n106;
  assign n108 = ~n80 & n107;
  assign n109 = ~n85 & n108;
  assign n110 = ~n90 & n109;
  assign n111 = ~n95 & n110;
  assign n112 = ~n100 & n111;
  assign 329 = n105 | ~n112;
  assign n114 = ~n65 & ~329;
  assign n115 = n65 & 329;
  assign n116 = ~n114 & ~n115;
  assign n117 = 4 & ~14;
  assign n118 = ~n63 & n117;
  assign n119 = ~n116 & n118;
  assign n120 = ~n70 & ~329;
  assign n121 = n70 & 329;
  assign n122 = ~n120 & ~n121;
  assign n123 = 17 & ~27;
  assign n124 = ~n68 & n123;
  assign n125 = ~n122 & n124;
  assign n126 = ~n75 & ~329;
  assign n127 = n75 & 329;
  assign n128 = ~n126 & ~n127;
  assign n129 = 30 & ~40;
  assign n130 = ~n73 & n129;
  assign n131 = ~n128 & n130;
  assign n132 = ~n80 & ~329;
  assign n133 = n80 & 329;
  assign n134 = ~n132 & ~n133;
  assign n135 = 43 & ~53;
  assign n136 = ~n78 & n135;
  assign n137 = ~n134 & n136;
  assign n138 = ~n85 & ~329;
  assign n139 = n85 & 329;
  assign n140 = ~n138 & ~n139;
  assign n141 = 56 & ~66;
  assign n142 = ~n83 & n141;
  assign n143 = ~n140 & n142;
  assign n144 = ~n90 & ~329;
  assign n145 = n90 & 329;
  assign n146 = ~n144 & ~n145;
  assign n147 = 69 & ~79;
  assign n148 = ~n88 & n147;
  assign n149 = ~n146 & n148;
  assign n150 = ~n95 & ~329;
  assign n151 = n95 & 329;
  assign n152 = ~n150 & ~n151;
  assign n153 = 82 & ~92;
  assign n154 = ~n93 & n153;
  assign n155 = ~n152 & n154;
  assign n156 = ~n100 & ~329;
  assign n157 = n100 & 329;
  assign n158 = ~n156 & ~n157;
  assign n159 = 95 & ~105;
  assign n160 = ~n98 & n159;
  assign n161 = ~n158 & n160;
  assign n162 = ~n105 & ~329;
  assign n163 = n105 & 329;
  assign n164 = ~n162 & ~n163;
  assign n165 = 108 & ~115;
  assign n166 = ~n103 & n165;
  assign n167 = ~n164 & n166;
  assign n168 = ~n119 & ~n125;
  assign n169 = ~n131 & n168;
  assign n170 = ~n137 & n169;
  assign n171 = ~n143 & n170;
  assign n172 = ~n149 & n171;
  assign n173 = ~n155 & n172;
  assign n174 = ~n161 & n173;
  assign 370 = n167 | ~n174;
  assign n176 = \1  & 223;
  assign n177 = 8 & 329;
  assign n178 = 14 & 370;
  assign n179 = 4 & ~n176;
  assign n180 = ~n177 & n179;
  assign n181 = ~n178 & n180;
  assign n182 = 11 & 223;
  assign n183 = 21 & 329;
  assign n184 = 27 & 370;
  assign n185 = ~n182 & ~n183;
  assign n186 = ~n184 & n185;
  assign n187 = 17 & n186;
  assign n188 = 24 & 223;
  assign n189 = 34 & 329;
  assign n190 = 40 & 370;
  assign n191 = ~n188 & ~n189;
  assign n192 = ~n190 & n191;
  assign n193 = 30 & n192;
  assign n194 = 37 & 223;
  assign n195 = 47 & 329;
  assign n196 = 53 & 370;
  assign n197 = ~n194 & ~n195;
  assign n198 = ~n196 & n197;
  assign n199 = 43 & n198;
  assign n200 = 50 & 223;
  assign n201 = 60 & 329;
  assign n202 = 66 & 370;
  assign n203 = ~n200 & ~n201;
  assign n204 = ~n202 & n203;
  assign n205 = 56 & n204;
  assign n206 = 63 & 223;
  assign n207 = 73 & 329;
  assign n208 = 79 & 370;
  assign n209 = ~n206 & ~n207;
  assign n210 = ~n208 & n209;
  assign n211 = 69 & n210;
  assign n212 = 76 & 223;
  assign n213 = 86 & 329;
  assign n214 = 92 & 370;
  assign n215 = ~n212 & ~n213;
  assign n216 = ~n214 & n215;
  assign n217 = 82 & n216;
  assign n218 = 89 & 223;
  assign n219 = 99 & 329;
  assign n220 = 105 & 370;
  assign n221 = ~n218 & ~n219;
  assign n222 = ~n220 & n221;
  assign n223 = 95 & n222;
  assign n224 = 102 & 223;
  assign n225 = 112 & 329;
  assign n226 = 115 & 370;
  assign n227 = ~n224 & ~n225;
  assign n228 = ~n226 & n227;
  assign n229 = 108 & n228;
  assign n230 = ~n187 & ~n193;
  assign n231 = ~n199 & n230;
  assign n232 = ~n205 & n231;
  assign n233 = ~n211 & n232;
  assign n234 = ~n217 & n233;
  assign n235 = ~n223 & n234;
  assign n236 = ~n229 & n235;
  assign 421 = ~n181 & ~n236;
  assign n238 = ~n193 & n199;
  assign n239 = n230 & ~n238;
  assign 430 = n205 | ~n239;
  assign n241 = ~n193 & ~n199;
  assign n242 = n211 & n241;
  assign n243 = ~n205 & n242;
  assign n244 = ~n199 & ~n205;
  assign n245 = n217 & n244;
  assign n246 = n230 & ~n243;
  assign 431 = n245 | ~n246;
  assign n248 = ~n217 & n241;
  assign n249 = n223 & n248;
  assign n250 = ~n187 & ~n238;
  assign n251 = ~n243 & n250;
  assign 432 = n249 | ~n251;
endmodule


