module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, y0, y1, y2, y3, y4);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10;
  output y0, y1, y2, y3, y4;
  wire n12, n13, n14, n15, n16, n17, n18, n19, n20, n21;
  assign n12 = x1 | x6;
  assign n13 = x0 & x4;
  assign n14 = x2 | n13;
  assign n15 = x3 | x5;
  assign n16 = (x3 & n14) | (x3 & n15) | (n14 & n15);
  assign n17 = (x1 & n12) | (x1 & n16) | (n12 & n16);
  assign n18 = x9 | x10;
  assign n19 = x7 | x8;
  assign n20 = (x7 & n17) | (x7 & n19) | (n17 & n19);
  assign n21 = (x10 & n18) | (x10 & n20) | (n18 & n20);
  assign y0 = n17;
  assign y1 = n16;
  assign y2 = n14;
  assign y3 = n21;
  assign y4 = n20;
endmodule
